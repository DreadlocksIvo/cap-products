ID,Description,ShortDescription
1,,