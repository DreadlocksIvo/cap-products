ID,DeliveryDate,Revenue
,,