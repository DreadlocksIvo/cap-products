ID,Description
BB,