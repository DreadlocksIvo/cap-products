ID,Name,Street,City,State,PostalCode,Country,Email,Phone,Fax
AA,,,,,,,,,