ID,Name
BB,