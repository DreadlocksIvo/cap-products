Name,Rating,Comment
,,