ID,Name,address_Street,address_City,address_State,address_PostalCode,address_Country,Email,Phone,Fax
AA,,,,,,,,,